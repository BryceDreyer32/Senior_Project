module temp (
    input clk,
    output o
);

assign o = clk;
endmodule
