module top();
/*angle_to_pwm a2p1(
    .reset_n,        // Active low reset
    .clock,          // The main clock
    .target_angle,   // The angle the wheel needs to move to in degrees. This number is multiplied by 2 internally
    .current_angle,  // The angle read from the motor encoder
    .pwm_done,       // Indicator from PWM that the pwm_ratio has been applied
    .angle_update,   // Request to update the angle
    .angle_done,     // Indicator that the angle has been applied 
    .pwm_update,     // Request an update to the PWM ratio
    .pwm_ratio,      // The high-time of the PWM signal out of 255.
    .pwm_direction   // The direction of the motor
);*/
endmodule